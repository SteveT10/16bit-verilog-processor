module Datapath();



endmodule